//PACKAGE

`include "apb_interface.sv"
package apb_pkg;

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "apb_master_transaction.sv"
`include "apb_slave_transcation.sv"
`include "apb_slave_config.sv"
`include "apb_master_sequencer.sv"
`include "apb_slave_sequencer.sv" 
`include "apb_master_driver.sv"
`include "apb_slave_driver.sv"
`include "apb_master_monitor.sv"
`include "apb_slave_monitor.sv"
`include "apb_master_sequence.sv"
`include "apb_slave_sequence.sv"  
 `include "apb_master_agent.sv"
 
`include "apb_slave_agent.sv"
`include "apb_env.sv"
`include "apb_test.sv"
`include "apb_high_range_pwdata.sv"
`include "apb_high_range_paddr.sv"
`include "apb_low_range_paddr.sv"
`include "apb_low_range_pwdata.sv"
`include "apb_test_high_range_pwdata.sv"
`include "apb_test_high_range_paddr.sv"
`include "apb_test_low_range_paddr.sv"
`include "apb_test_low_range_pwdata.sv"


endpackage
 
 
 
 
  



